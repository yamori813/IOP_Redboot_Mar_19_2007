# ====================================================================
#
#      hal_arm_xscale_iop33x.cdl
#
#      Intel XScale architectural HAL package configuration data
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 1998, 1999, 2000, 2001, 2002, 2003 Red Hat, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
## at http://sources.redhat.com/ecos/ecos-license/
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      drew.moseley@intel.com
# Original data:  msalter
# Contributors:
# Date:           2003-07-10
#
# Copyright:    (C) 2003-2004 Intel Corporation.
#####DESCRIPTIONEND####
#
# ====================================================================
cdl_package CYGPKG_HAL_ARM_XSCALE_IOP33X {
    display       "Intel XScale IOP331 and IOP332 IO Processors"
    parent        CYGPKG_HAL_ARM_XSCALE_IOP
    hardware
    include_dir   cyg/hal
    define_header hal_arm_xscale_iop33x.h
    requires      CYGSEM_HAL_ARM_XSCALE_IOP_PROVIDE_I2C_API
    requires      { !CYGPKG_REDBOOT || CYGSEM_HAL_ARM_XSCALE_IOP_PROVIDE_PCI_REDBOOT_FNS }
    requires      { !CYGPKG_REDBOOT || CYGSEM_HAL_ARM_XSCALE_IOP_PROVIDE_ECC_REDBOOT_FNS }
    requires      { CYGNUM_HAL_ARM_XSCALE_IOP_NUM_BARS == 4 }
    description   "
        This HAL variant package provides generic
        support for the Intel IOP331 and IOP332 IO processors.
        It is also necessary to select a specific target platform
        HAL package."

    # Let the architectural HAL see this variant's interrupts file
     define_proc {
        puts $::cdl_header \
       "#define CYGBLD_HAL_VAR_INTS_H <cyg/hal/hal_var_ints.h>"
        puts $::cdl_header \
       "#define CYGBLD_HAL_VAR_H <cyg/hal/hal_iop33x.h>"

        puts $::cdl_system_header "#define CYGBLD_HAL_ARM_VAR_IO_H"
    }

    compile       iop33x_misc.c iop33x_pci.c

    # Real-time clock/counter specifics
    cdl_component CYGNUM_HAL_RTC_CONSTANTS {
        display       "Real-time clock constants"
        flavor        none
        no_define
    
        cdl_option CYGNUM_HAL_RTC_NUMERATOR {
            display       "Real-time clock numerator"
            flavor        data
            calculated    1000000000
        }
        cdl_option CYGNUM_HAL_RTC_DENOMINATOR {
            display       "Real-time clock denominator"
            flavor        data
            default_value 100
            description   "
              This option selects the heartbeat rate for the real-time clock.
              The rate is specified in ticks per second.  Change this value
              with caution - too high and your system will become saturated
              just handling clock interrupts, too low and some operations
              such as thread scheduling may become sluggish."
        }
        cdl_option CYGNUM_HAL_RTC_PERIOD {
            display       "Real-time clock period"
            flavor        data
            calculated    1000000/CYGNUM_HAL_RTC_DENOMINATOR
	    description   "
              This value gives the RTC period in microseconds. It is
              translated into the actual clock period value in the clock
              init and read functions."
        }
    }

    # ECC Memory Configuration
    cdl_component CYGNUM_HAL_ECC_CONFIGURATION {
        display       "ECC Memory Configuration"
        flavor        none
        no_define

        cdl_option CYGSEM_HAL_ARM_IOP33X_ENABLE_ECC {
            display       "Enable ECC region"
            flavor        bool
            default_value 1
            description   "
            This option controls whether or not the HAL will enable ECC."
        }

        cdl_option CYGSEM_HAL_ARM_IOP33X_32BIT_ECC_REGION_SIZE {
            display       "Enable 32-bit ECC region of a given size in megabytes"
            flavor        data
            default_value { (CYGSEM_HAL_ARM_IOP33X_ENABLE_ECC == 1) ? 0 : 0 }
            active_if     { CYGSEM_HAL_ARM_IOP33X_ENABLE_ECC == 1 }
            legal_values  0 1 2 4 8 16 32 64 128 256 512
            description   "
            This option controls the size of the 32-bit ECC region."
        }
    }

    cdl_component CYGPKG_REDBOOT_XSCALE_OPTIONS {
        display       "Redboot for XScale options"
        flavor        none
        no_define
        parent        CYGPKG_REDBOOT
        active_if     CYGPKG_REDBOOT
        description   "
            This option lists the target's requirements for a valid Redboot
            configuration."

        # RedBoot details
        requires { !CYGPKG_REDBOOT_ARM_LINUX_EXEC || \
                       CYGHWR_REDBOOT_ARM_LINUX_EXEC_ADDRESS_DEFAULT == 0xA0008000 }
        define_proc {
            puts $::cdl_header "#define CYGHWR_REDBOOT_ARM_TRAMPOLINE_ADDRESS 0x00001f00"
        }
    }

    cdl_component CYGPKG_REDBOOT_PLATFORM_MEMORY_INFO {
        display       "Print platform-specific memory information"
        flavor        none
        no_define
        parent        CYGPKG_REDBOOT
        active_if     CYGPKG_REDBOOT
        description   "
            This option enables platform-specific memory information to be printed."

        define_proc {
            puts $::cdl_header "#define HAL_PLATFORM_MEMORY_INFO hal_platform_memory_info"
        }
    }
}
