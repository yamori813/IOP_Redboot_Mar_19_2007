# ====================================================================
#
#      hal_arm_xscale_core.cdl
#
#      Intel XScale architectural HAL package configuration data
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 1998, 1999, 2000, 2001, 2002, 2003, 2004 Red Hat, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
## at http://sources.redhat.com/ecos/ecos-license/
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      msalter
# Original data:  msalter, dmoseley, cbruns
# Contributors:
# Date:           2002-10-18
#
# Copyright:    (C) 2003-2004 Intel Corporation.
#####DESCRIPTIONEND####
#
# ====================================================================
cdl_package CYGPKG_HAL_ARM_XSCALE_CORE {
    display       "Intel XScale Core Support"
    parent        CYGPKG_HAL_ARM
    hardware
    include_dir   cyg/hal
    define_header hal_arm_xscale_core.h
    description   "
        This HAL variant package provides generic support common
        to Intel XScale CPU cores. It is also necessary to select
        a specific target platform and CPU HAL package."

    implements    CYGINT_HAL_ARM_ARCH_XSCALE

    compile       xscale_misc.c xscale_stub.c

    cdl_option CYGSEM_HAL_ARM_XSCALE_BTB {
    	display       "Enable Branch Target Buffer"
        flavor        bool
        default_value 1
        description   "
            This option controls whether or not the Branch Target
            Buffer is enabled. The BTB is used for branch prediction
            and can have significant performance benefits. Control
            is provided because there is an errata for A-step 80200
            CPUS which will lead to problems with thumb branches
            if the BTB is on. Normal ARM programs are not affected
            by this errata."
    }

    cdl_option CYGSEM_HAL_ARM_XSCALE_USE_CACHE_AS_SRAM {
        display "Lock the DCache at base of RAM"
        flavor  bool
        default_value 0
        # Currently only implemented on the IQ80331/IQ80332 and IQ8134X CRBs
        requires { CYGPKG_HAL_ARM_XSCALE_IQ8033X || CYGPKG_HAL_ARM_XSCALE_IQ8134X }
        requires CYGSEM_HAL_BUILD_MINIMAL_REDBOOT
        requires { CYG_HAL_STARTUP=="ROM" }
        requires { CYG_HAL_STARTUP_EXTRA=="-CACHE-SRAM" }
        description   "
                This option controls whether the HAL will lock the DCache at the base
                of RAM.  This allows the DCache to be effectively used as SRAM and
                will allow a certain amount of functionality even if no SDRAM is
                present."
    }

    cdl_option CYGSEM_HAL_ARM_HOTDEBUG {
            display       "Add Hot Debug support"
            flavor        bool
            default_value 0
            description   "
                This option adds in JTAG Hot Debug support code to the
                RESET vector start up code. _xscale_hotdebug... Macros
                are located in hal_hotdebug.h "
        }
 cdl_option CYGNUM_HAL_ARM_XSCALE_CORE_GENERATION {
        display       "XScale core generation"
        flavor        data
        legal_values  1 2 3 
        default_value 1
        description   "
            This option selects the XScale generation for the core
            being used in a particular IOP."
    }

    cdl_option CYGNUM_HAL_ARM_XSCALE_IOP_GENERATION {
        display       "IOP generation"
        flavor        data
        legal_values  1 2 3 4 
        default_value 1
        description   "
            This option selects the IOP generation."
	}
	cdl_option CYGSEM_HAL_ENABLE_L2_CACHE {
        display       "Enable L2 Cache"
        active_if { (CYGNUM_HAL_ARM_XSCALE_CORE_GENERATION > 2)  } 
        flavor        bool 
        default_value 1
        description   "
            Select whether or not the L2 Cache should be enabled."
    }
}
