# ====================================================================
#
#      hal_arm_xscale_iq80315.cdl
#
#      Intel XScale IQ80315 platform HAL package configuration data
#
# ====================================================================
#####COPYRIGHTBEGIN####
#
# -------------------------------------------
# The contents of this file are subject to the Red Hat eCos Public License
# Version 1.1 (the "License"); you may not use this file except in
# compliance with the License.  You may obtain a copy of the License at
# http://www.redhat.com/
#
# Software distributed under the License is distributed on an "AS IS"
# basis, WITHOUT WARRANTY OF ANY KIND, either express or implied.  See the
# License for the specific language governing rights and limitations under
# the License.
#
# The Original Code is eCos - Embedded Configurable Operating System,
# released September 30, 1998.
#
# The Initial Developer of the Original Code is Red Hat.
# Portions created by Red Hat are
# Copyright (C) 1998, 1999, 2000, 2001 Red Hat, Inc.
# All Rights Reserved.
# -------------------------------------------
#
#####COPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      dkranak
# Contributors:   hmt
# Date:           2001-12-03
#
# Copyright:    (C) 2003-2004 Intel Corporation.
#####DESCRIPTIONEND####
#
# ====================================================================
cdl_package CYGPKG_HAL_ARM_XSCALE_IQ80315 {
    display       "Intel XScale IQ80315 evaluation board"
    parent        CYGPKG_HAL_ARM_XSCALE
    hardware
    include_dir   cyg/hal
    define_header hal_arm_xscale_iq80315.h
    description   "
        This HAL platform package provides
        support for the Intel XScale IQ80315 board."

    compile       iq80315_misc.c iq80315_pci.c iq80315_cf.c

    implements    CYGINT_HAL_DEBUG_GDB_STUBS
    implements    CYGINT_HAL_DEBUG_GDB_STUBS_BREAK
    implements    CYGINT_HAL_VIRTUAL_VECTOR_SUPPORT
    implements    CYGINT_HAL_ARM_MEM_REAL_REGION_TOP
    implements    CYGINT_HAL_VIRTUAL_VECTOR_COMM_BAUD_SUPPORT

    include_dir    cyg/hal

    define_proc {
        puts $::cdl_system_header "#define CYGBLD_HAL_TARGET_H   <pkgconf/hal_arm.h>"
        puts $::cdl_system_header "#define CYGBLD_HAL_VARIANT_H  <pkgconf/hal_arm_xscale_ioc80314.h>"
        puts $::cdl_system_header "#define CYGBLD_HAL_PLATFORM_H <pkgconf/hal_arm_xscale_iq80315.h>"
        puts $::cdl_system_header "#define CYGBLD_HAL_BOARD_H    <cyg/hal/iq80315.h>"
        puts $::cdl_system_header "#define CYGBLD_HAL_DIAG_INL   <cyg/hal/hal_diag_iq80315.inl>"
        puts $::cdl_header "#define CYGBLD_HAL_PLF_INTS_H <cyg/hal/hal_plf_ints.h>"
	puts $::cdl_header "#define HAL_PLATFORM_CPU    \"XScale\""
        puts $::cdl_header "#define HAL_PLATFORM_MACHINE_TYPE  353"
# This is defined in iq80315.h        puts $::cdl_header "#define HAL_PLATFORM_BOARD  \"IQ80315\""
# This is defined in iq80315.h       puts $::cdl_header "#define HAL_PLATFORM_EXTRA  \"\""
    }

    cdl_component CYG_HAL_STARTUP {
        display       "Startup type"
        flavor        data
        default_value {"RAM"}
        legal_values  {"RAM" "ROM"}
	no_define
	define -file system.h CYG_HAL_STARTUP
        description   "
           When targeting the IQ80315 eval board it is possible to build
           the system for either RAM bootstrap or ROM bootstrap(s). Select
           'ram' when building programs to load into RAM using onboard
           debug software such as Angel or eCos GDB stubs.  Select 'rom'
           when building a stand-alone application which will be put
           into ROM.  Selection of 'stubs' is for the special case of
           building the eCos GDB stubs themselves."
    }

        cdl_option NUM_HAL_CPU_0_BASE_PHY_ADDR {
            display       "CPU 0 base physical address."
            flavor        data
            default_value 0x00000000
            define -file system.h NUM_HAL_CPU_0_BASE_PHY_ADDR
            description   "
                Defines CPU 0 physical varialble address space."
        }

        cdl_option NUM_HAL_CPU_0_BASE_VIR_ADDR {
            display       "CPU 0 base virtural address."
            flavor        data
            default_value 0x00000000
            define -file system.h NUM_HAL_CPU_0_BASE_VIR_ADDR
            description   "
                Defines CPU 0 virtural varialble address space."
        }

        cdl_option NUM_HAL_CPU_0_VAR_SIZE {
            display       "CPU 0 base virtural address size."
            flavor        data
            default_value 0x00100000
            define -file system.h NUM_HAL_CPU_0_VAR_SIZE
            description   "
                Defines size of CPU 0 varialble address space."
        }

    cdl_component PKG_HAL_HAS_MULT_CPU {
        display "Intel XScale IQ80315 Supports Muliplal Processors"
            default_value 1
        description   "
            Package specific support for more than one processor."

        cdl_option NUM_HAL_CPU_1_BASE_PHY_ADDR {
            display       "CPU 1 base physical address."
            flavor        data
            default_value 0x00100000
            define -file system.h NUM_HAL_CPU_1_BASE_PHY_ADDR
            description   "
                Defines CPU 1 physical variable address space."
        }

        cdl_option NUM_HAL_CPU_1_BASE_VIR_ADDR {
            display       "CPU 1 base virtural address."
            flavor        data
            default_value 0x00000000
            define -file system.h NUM_HAL_CPU_0_BASE_VIR_ADDR
            description   "
                Defines CPU 1 virtural varialble address space."
        }

        cdl_option NUM_HAL_CPU_1_VAR_SIZE {
            display       "CPU 1 base virtural address size."
            flavor        data
            default_value 0x00100000
            define -file system.h NUM_HAL_CPU_1_VAR_SIZE
            description   "
                Defines size of CPU 1 varialble address space."
        }


    }

    cdl_component CYGPKG_HAL_ARM_XSCALE_IQ80315_COMPONENT_SETTINGS {
        display "Intel XScale IQ80315 Component Settings"
        flavor  none
        no_define
        description   "
            Package specific component base address and initial
            values."

        cdl_option HAL_IOC80314_CSR_BASE {
            display       "Relocated base address of CSR Reg."
            flavor        data
            default_value 0x50100000
            define -file system.h HAL_IOC80314_CSR_BASE
            description   "
                Relocated base address of Control Space Registes.  The default value
                after Reset is 0xFFFE0000.  This value is placed into CIU_CFG_BAR at
                the beginning of the processor boot code."
        }

        cdl_option HAL_IOC80314_SDRAM_VIR_BASE {
            display       "SDRAM Virtual Base address."
            flavor        data
            default_value 0x00000000
            define -file system.h HAL_IOC80314_SDRAM_VIR_BASE
            description   "
                Defines base address of SDRAM (virtual)."
        }

        cdl_option HAL_IOC80314_FLASH_BASE {
            display       "Relocated FLASH base address."
            flavor        data
            default_value 0x40000000
            define -file system.h HAL_IOC80314_FLASH_BASE
            description   "
                Relocated FLASH base address attached to signal PCE0#.  The default value
                after Reset is 0x00000000.  This value is placed into CIU_SF_BAR1 at
                the beginning of the processor boot code."
        }

        cdl_option HAL_IOC80314_SRAM_BASE {
            display       "Relocated FLASH base address."
            flavor        data
            default_value 0x50000000
            define -file system.h HAL_IOC80314_SRAM_BASE
            description   "
                SRAM base address location.  The default value
                after Reset is undefined and disabled.  This value is placed into
                CIU_SRAM_BAR at the beginning of the processor boot code."
        }

        cdl_option HAL_IOC80314_SRAM_SIZE {
            display       "Size size."
            flavor        data
            legal_values  {0x0 0x100000}
            default_value 0x100000
            define -file system.h HAL_IOC80314_SRAM_SIZE
            description   "
                SRAM size in bytes."
        }
        cdl_option HAL_IOC80314_CIU_PCI1_BASE {
            display       "CIU base address to access PCI1."
            flavor        data
            default_value 0x80000000
            define -file system.h HAL_IOC80314_CIU_PCI1_BASE
            description   "
                CIU base address location to access PCI1 through the SFN.  The default value
                after Reset is undefined and disabled.  This value is placed into
                CIU_BAR2 at PCI init."
        }

        cdl_option HAL_IOC80314_CIU_PCI2_BASE {
            display       "CIU base address to access PCI1."
            flavor        data
            default_value 0xC0000000
            define -file system.h HAL_IOC80314_CIU_PCI2_BASE
            description   "
                CIU base address location to access PCI1 through the SFN.  The default value
                after Reset is undefined and disabled.  This value is placed into
                CIU_BAR2 at PCI init."
        }
    }

    cdl_option CYGNUM_HAL_PROCESSOR_SPEED {
        display       "Clock speed of the processor"
        flavor        data
        legal_values  5000000 100000000
        default_value 100000000;
        description   "
            This option selects the operating frequency of the processor."
    }

    cdl_option CYGNUM_HAL_SFN_SPEED {
        display       "ioc80314 SFN speed"
        flavor        data
        legal_values  5000000 133000000 100000000
        default_value 133000000;
        description   "
            This option selects the operating frequency of the
            ioc80314 internal Switch Fabric Network.  This is used
            to define the UART clock speed and PBI interface timings."
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL_BAUD {
        display       "Diagnostic serial port baud rate"
        flavor        data
        legal_values  9600 19200 38400 57600 115200
        default_value 115200   ;
        description   "
            This option selects the baud rate used for the diagnostic port.
            Note: this should match the value chosen for the GDB port if the
            diagnostic and GDB port are the same."
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL_BAUD {
        display       "GDB serial port baud rate"
        flavor        data
        legal_values  9600 19200 38400 57600 115200
        default_value 115200   ;
        description   "
            This option selects the baud rate used for the diagnostic port.
            Note: this should match the value chosen for the GDB port if the
            diagnostic and GDB port are the same."
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS {
        display      "Number of communication channels on the board"
        flavor       data
        calculated   2
	description "
	    Channel 0 is the only serial port on the board."
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL {
        display          "Debug serial port"
        active_if        CYGPRI_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL_CONFIGURABLE
        flavor data
        legal_values     0 to CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS-1
        default_value    0
        description      "
            The IQ80315 has only one serial port."
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL {
	display          "Diagnostic serial port"
        active_if        CYGPRI_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL_CONFIGURABLE
	flavor data
	legal_values     0 to CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS-1
	default_value    0
	description      "
            The IQ80315 has only one serial port."
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL_DEFAULT {
        display      "Default console channel."
        flavor       data
        legal_values     0 to CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS-1
        calculated   0
    }

    cdl_component CYGBLD_GLOBAL_OPTIONS {
        display "Global build options"
        flavor  none
        no_define
        description   "
	    Global build options including control over
	    compiler flags, linker flags and choice of toolchain."

        parent  CYGPKG_NONE

        cdl_option CYGBLD_GLOBAL_COMMAND_PREFIX {
            display "Global command prefix"
            flavor  data
            no_define
            default_value { "xscale-elf" }
            description "
                This option specifies the command prefix used when
                invoking the build tools."
        }

        cdl_option CYGBLD_GLOBAL_CFLAGS {
            display "Global compiler flags"
            flavor  data
            no_define
            default_value { "-mcpu=xscale -Wall -Wpointer-arith -Wstrict-prototypes -Winline -Wundef -Woverloaded-virtual -g -O2 -ffunction-sections -fdata-sections -fno-rtti -fno-exceptions -fvtable-gc -finit-priority -mapcs-frame" }
            description   "
                This option controls the global compiler flags which are used to
                compile all packages by default. Individual packages may define
                options which override these global flags."
        }

        cdl_option CYGBLD_GLOBAL_LDFLAGS {
            display "Global linker flags"
            flavor  data
            no_define
            ###default_value { "-mcpu=xscale -Wl,--gc-sections -Wl,-static -g -O2 -nostdlib -Wl,--cref,-Map,$(PREFIX)/bin/redboot.map -Wl,--verbose" }
            default_value { "-mcpu=xscale -Wl,--gc-sections -Wl,-static -g -O2 -nostdlib -Wl,--cref,-Map,$(PREFIX)/bin/redboot.map" }
            description   "
                This option controls the global linker flags. Individual
                packages may define options which override these global flags."
        }

        cdl_option CYGBLD_BUILD_GDB_STUBS {
            display "Build GDB stub ROM image"
            default_value 0
            requires { CYG_HAL_STARTUP == "ROM" }
            requires CYGSEM_HAL_ROM_MONITOR
            requires CYGBLD_BUILD_COMMON_GDB_STUBS
            requires CYGDBG_HAL_DEBUG_GDB_INCLUDE_STUBS
            requires CYGDBG_HAL_DEBUG_GDB_BREAK_SUPPORT
            requires CYGDBG_HAL_DEBUG_GDB_THREAD_SUPPORT
            requires ! CYGDBG_HAL_COMMON_INTERRUPTS_SAVE_MINIMUM_CONTEXT
            requires ! CYGDBG_HAL_COMMON_CONTEXT_SAVE_MINIMUM
            no_define
            description "
                This option enables the building of the GDB stubs for the
                board. The common HAL controls takes care of most of the
                build process, but the final conversion from ELF image to
                binary data is handled by the platform CDL, allowing
                relocation of the data if necessary."

            make -priority 320 {
                <PREFIX>/bin/gdb_module.bin : <PREFIX>/bin/gdb_module.img
                $(OBJCOPY) --remove-section=.fixed_vectors -O binary $< $@
            }
        }
    }

    cdl_component CYGPKG_HAL_ARM_XSCALE_IQ80315_OPTIONS {
        display "Intel XScale IQ80315 build options"
        flavor  none
        no_define
        description   "
	    Package specific build options including control over
	    compiler flags used only in building this package,
	    and details of which tests are built."

        cdl_option CYGPKG_HAL_ARM_XSCALE_IQ80315_BOARD_FLAVOR {
            display "Different Options for different Flavors"
            flavor  data
	    default_value {"IQ80315"}
	    legal_values  {"IQ80315" "XCARD"}
	    define -file system.h CYGPKG_HAL_ARM_XSCALE_IQ80315_BOARD_FLAVOR
            description   "
                This option will change some settings based on the board flavor."
		
        }

        cdl_option CYGPKG_HAL_ARM_XSCALE_IQ80315_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the XScale IQ80315 HAL. These flags are used in addition
                to the set of global flags."
        }

        cdl_option CYGPKG_HAL_ARM_XSCALE_IQ80315_CFLAGS_REMOVE {
            display "Suppressed compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the XScale IQ80315 HAL. These flags are removed from
                the set of global flags if present."
        }

	cdl_option CYGNUM_HAL_BREAKPOINT_LIST_SIZE {
            display       "Number of breakpoints supported by the HAL."
            flavor        data
            default_value 32
            description   "
                This option determines the number of breakpoints supported by the HAL."
        }
    }

    cdl_component CYGHWR_MEMORY_LAYOUT {
        display "Memory layout"
        flavor data
        no_define
        calculated { CYG_HAL_STARTUP == "RAM" ? "arm_xscale_iq80315_ram" : \
                                                "arm_xscale_iq80315_rom" }

        cdl_option CYGHWR_MEMORY_LAYOUT_LDI {
            display "Memory layout linker script fragment"
            flavor data
            no_define
            define -file system.h CYGHWR_MEMORY_LAYOUT_LDI
            calculated { CYG_HAL_STARTUP == "RAM" ? "<pkgconf/mlt_arm_xscale_iq80315_ram.ldi>" : \
                                                    "<pkgconf/mlt_arm_xscale_iq80315_rom.ldi>" }
        }

        cdl_option CYGHWR_MEMORY_LAYOUT_H {
            display "Memory layout header file"
            flavor data
            no_define
            define -file system.h CYGHWR_MEMORY_LAYOUT_H
            calculated { CYG_HAL_STARTUP == "RAM" ? "<pkgconf/mlt_arm_xscale_iq80315_ram.h>" : \
                                                    "<pkgconf/mlt_arm_xscale_iq80315_rom.h>" }
        }
    }

    cdl_option CYGSEM_HAL_ROM_MONITOR {
        display       "Behave as a ROM monitor"
        flavor        bool
        default_value 0
        parent        CYGPKG_HAL_ROM_MONITOR
        requires      { CYG_HAL_STARTUP == "ROM" }
        description   "
            Enable this option if this program is to be used as a ROM monitor,
            i.e. applications will be loaded into RAM on the board, and this
            ROM monitor may process exceptions or interrupts generated from the
            application. This enables features such as utilizing a separate
            interrupt stack when exceptions are generated."
    }

    cdl_option CYGSEM_HAL_USE_ROM_MONITOR {
         display       "Work with a ROM monitor"
         flavor        booldata
         legal_values  { "Generic" "GDB_stubs" }
         default_value { CYG_HAL_STARTUP == "RAM" ? "GDB_stubs" : 0 }
         parent        CYGPKG_HAL_ROM_MONITOR
         requires      { CYG_HAL_STARTUP == "RAM" }
         description   "
             Support can be enabled for different varieties of ROM monitor.
             This support changes various eCos semantics such as the encoding
             of diagnostic output, or the overriding of hardware interrupt
             vectors.
             Firstly there is \"Generic\" support which prevents the HAL
             from overriding the hardware vectors that it does not use, to
             instead allow an installed ROM monitor to handle them. This is
             the most basic support which is likely to be common to most
             implementations of ROM monitor.
             \"GDB_stubs\" provides support when GDB stubs are included in
             the ROM monitor or boot ROM."
     }

    cdl_component CYGPKG_REDBOOT_HAL_OPTIONS {
        display       "Redboot HAL options"
        flavor        none
        no_define
        parent        CYGPKG_REDBOOT
        active_if     CYGPKG_REDBOOT
        description   "
            This option lists the target's requirements for a valid Redboot
            configuration."

        # compile -library=libextras.a redboot_cmds.c

        cdl_option CYGBLD_BUILD_REDBOOT_BIN {
            display       "Build Redboot ROM binary image"
            active_if     CYGBLD_BUILD_REDBOOT
            default_value 1
            no_define
            description "This option enables the conversion of the Redboot ELF
                         image to a binary image suitable for ROM programming."

            compile -library=libextras.a                                   \
                                diag/diag.c                                \
                                diag/io_utils.c                            \
                                diag/xscale_test.c                         \
                                diag/memtest.c                             \
                                diag/test_menu.c                           \
                                diag/bootE2.c                              \
                                diag/pcitest.c                             \
                                diag/battery.c                             \
                                diag/lcd.c                                 \
                                diag/timer.c                               \
                                diag/rtc.c                                 \
                                diag/cftest.c                              \
                                diag/sata.c


            make -priority 325 {
                <PREFIX>/bin/redboot.bin : <PREFIX>/bin/redboot.elf
                $(OBJCOPY) --strip-debug $< $(@:.bin=.img)
                $(OBJCOPY) -O srec $< $(@:.bin=.srec)
                $(OBJCOPY) -O binary $< $@
            }
        }

        cdl_option CYGSEM_HAL_ARM_IQ80315_BATTERY_TEST {
            display       "Include Battery Test in Diagnostics Menu"
            flavor        bool
            default_value 1
            description   "
                This option controls whether or not the battery test is included
                in the IQ80315 diagnostics."
        }

        cdl_option CYGSEM_HAL_ROM_RESET_USES_JUMP {
            display       "Enables branch at reset instruction vector."
            flavor        bool
            default_value 1
            description   "
                This allows a branch instructon at address 0x00000000 thus
                provideing a position independent code for the reset
                instruction vector."
        }

    }

}
