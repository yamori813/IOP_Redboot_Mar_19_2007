# ====================================================================
#
#	intel_ioc80314_eth_drivers.cdl
#
#	Intel IOC80314 ethernet driver
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Red Hat, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
## at http://sources.redhat.com/ecos/ecos-license/
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      nickg, from i82559 original
# Original data:  hmt
# Contributors:	  hmt, gthomas, jskov, dkranak
# Date:           2001-10-25
# Copyright:    (C) 2003-2004 Intel Corporation.
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_DEVS_ETH_INTEL_IOC80314 {
    display       "Intel IOC80314 gigabit ethernet driver"
    description   "Ethernet driver for Intel IOC80314 Gigabit controller."

    parent        CYGPKG_IO_ETH_DRIVERS
    active_if     CYGPKG_IO_ETH_DRIVERS

    active_if     CYGINT_DEVS_ETH_INTEL_IOC80314_REQUIRED

    include_dir   cyg/devs/eth

    # SNMP demands to know stuff; this sadly makes us break the neat
    # abstraction of the device having nothing exported.
    include_files include/ioc80314_info.h SpacEthDefs.h SpacEthPublic.h SpacEthHardwareDefs.h tuntypes.h \
                   SpacRedBoot.h SpacQMng.h SpacEthRegOps.h	SpacEthInterrupts.h	\
				   SpacEthBuffDescript.h SpacEthArbitration.h 80200.h SpacSynch.h sys_utils.h ts_basic_types.h\
				   SpacEthDma.h	 SpacEthMac.h SpacEthMii.h

    # and tell them that it is available
    define_proc {
        puts $::cdl_header "#include CYGDAT_DEVS_ETH_INTEL_IOC80314_CFG";
    }

    compile       -library=libextras.a if_ioc80314.c SpacQMng.c SpacRedBoot.c SpacEthMii.c SpacEthDrv.c \
                           SpacEthRegOps.c sys_utils.c SpacEthArbitration.c  SpacEthInfo.c	 \
						   SpacEthMac.c	SpacEthBuffDescript.c SpacEthDma.c

    cdl_option CYGDBG_DEVS_ETH_INTEL_IOC80314_CHATTER {
	display "Prints ethernet device status info during startup"
        default_value 0
	description   "
	    The ethernet device initialization code can print lots of info
	    to confirm that it has found the devices on the PCI bus, read
	    the MAC address from EEPROM correctly, and so on
		"
    }

    cdl_option CYGDBG_DEVS_ETH_INTEL_IOC80314_INTERRUPT_DEBUG {
	display "Prints ethernet device status around interrupt routines"
	default_value 1
	description   "
	    The ethernet device initialization code can print info around
		the interrupt routines to assist in debugging.
		"
    }

    cdl_option CYGNUM_DEVS_ETH_INTEL_IOC80314_DEV_COUNT {
	display "Number of supported interfaces."
	calculated    { CYGINT_DEVS_ETH_INTEL_IOC80314_REQUIRED }
        flavor        data
	description   "
	    This option selects the number of gigE ports on the board
		"
    }

    cdl_component CYGDBG_DEVS_ETH_INTEL_IOC80314_KEEP_STATISTICS {
	display "Keep Ethernet statistics"
	default_value 0
	description   "
	    The ethernet device can maintain statistics about the network,
	    specifically a great variety of error rates which are useful
	    for network management.  SNMP for example uses this
	    information.  There is some performance cost in maintaining
	    this information; disable this option to recoup that."

	cdl_option CYGDBG_DEVS_ETH_INTEL_IOC80314_KEEP_IOC80314_STATISTICS {
	    display "Keep ioc80314 Internal statistics"
	    default_value 1
	    description   "
	        The ioc80314 keeps internal counters, and it is possible to
	        acquire these.  But the ioc80314 (reputedly) does not service
	        the network whilst uploading the data to RAM from its
	        internal registers.  If throughput is a problem, disable
	        this option to acquire only those statistics gathered by
	        software, so that the ioc80314 never sleeps."
	}
    }

    cdl_component CYGPKG_DEVS_ETH_INTEL_IOC80314_OPTIONS {
        display "Intel IOC80314 ethernet driver build options"
        flavor  none
	no_define

        cdl_option CYGPKG_DEVS_ETH_INTEL_IOC80314_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "-D_KERNEL -D__ECOS" }
            description   "
                This option modifies the set of compiler flags for
                building the Intel IOC80314 ethernet driver
                package. These flags are used in addition to the set of
                global flags."
        }
    }
}
# EOF intel_ioc80314_eth_drivers.cdl
